// Interfaces

module if2d
(
	input	clk,
	input	[1:0]	pattern,	//4x4, 8x8, 16x16
	
	output	res
);

assign res = clk;




endmodule

