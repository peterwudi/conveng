module ALU
(
	input		clk,
	
	output	res

);

assign res = clk;



endmodule

